`define AHB_HTRANS_IDLE 2'b00
`define AHB_HTRANS_BUSY 2'b01
`define AHB_HTRANS_NONSEQ 2'b10
`define AHB_HTRANS_SEQ 2'b11

`define AHB_HSIZE_BYTE 3'b000
`define AHB_HSIZE_HALFWORD 3'b001
`define AHB_HSIZE_WORD 3'b010
`define AHB_HSIZE_DOUBLEWORD 3'b011
`define AHB_HSIZE_4WORD 3'b100
`define AHB_HSIZE_8WORD 3'b101

`define AHB_HBURST_SINGLE 3'b000
`define AHB_HBURST_INCR 3'b001
`define AHB_HBURST_WRAP4 3'b010
`define AHB_HBURST_INCR4 3'b011
`define AHB_HBURST_WRAP8 3'b100
`define AHB_HBURST_INCR8 3'b101
`define AHB_HBURST_WRAP16 3'b110
`define AHB_HBURST_INCR16 3'b111

`define AHB_HRESP_OKAY 1'b0
`define AHB_HRESP_ERROR 1'b1

`define AVL_RESPONSE_OKAY 2'b00
`define AVL_RESPONSE_RESERVED 2'b01
`define AVL_RESPONSE_SLAVEERROR 2'b10
`define AVL_RESPONSE_DECODEERROR 2'b11
